module instr_mem (
    input logic clk,
    input logic [31:0] addr,
    output logic [31:0] instr
);
endmodule
