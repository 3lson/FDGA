// gpu_pynq_top.sv
`default_nettype none
`timescale 1ns/1ns

`include "common.svh"
`include "gpu_defines.svh" // Include your memory map defines

module gpu_pynq_top #(
    // Parameters for AXI Lite Interface
    parameter int C_S_AXI_DATA_WIDTH = 32,
    parameter int C_S_AXI_ADDR_WIDTH = 5, // 2^5 = 32 addresses for control

    // GPU Parameters
    parameter int DATA_MEM_NUM_CHANNELS      = 8,
    parameter int INSTRUCTION_MEM_NUM_CHANNELS = 8,
    parameter int NUM_CORES                  = 1,
    parameter int WARPS_PER_CORE             = 1,
    parameter int THREADS_PER_WARP           = 16
) (
    // AXI Lite Slave Interface (for PS control)
    input  wire                                 S_AXI_ACLK,
    input  wire                                 S_AXI_ARESETN,
    // ... standard AXI signals (AWADDR, WDATA, etc.). Vivado will connect these.
    input  wire [C_S_AXI_ADDR_WIDTH-1:0]        S_AXI_AWADDR,
    input  wire                                 S_AXI_AWVALID,
    output wire                                 S_AXI_AWREADY,
    input  wire [C_S_AXI_DATA_WIDTH-1:0]        S_AXI_WDATA,
    input  wire [C_S_AXI_DATA_WIDTH/8-1:0]      S_AXI_WSTRB,
    input  wire                                 S_AXI_WVALID,
    output wire                                 S_AXI_WREADY,
    output wire [1:0]                           S_AXI_BRESP,
    output wire                                 S_AXI_BVALID,
    input  wire                                 S_AXI_BREADY,
    input  wire [C_S_AXI_ADDR_WIDTH-1:0]        S_AXI_ARADDR,
    input  wire                                 S_AXI_ARVALID,
    output wire                                 S_AXI_ARREADY,
    output wire [C_S_AXI_DATA_WIDTH-1:0]        S_AXI_RDATA,
    output wire [1:0]                           S_AXI_RRESP,
    output wire                                 S_AXI_RVALID,
    input  wire                                 S_AXI_RREADY,

    // Instruction BRAM Interface
    output logic                                instr_bram_en,
    output logic [`INSTRUCTION_MEMORY_ADDRESS_WIDTH-1:0] instr_bram_addr,
    input  wire [`INSTRUCTION_WIDTH-1:0]        instr_bram_dout,

    // Data BRAM Interface
    output logic                                data_bram_en,
    output logic [`DATA_MEMORY_ADDRESS_WIDTH-1:0] data_bram_addr,
    output logic [0:0]                          data_bram_we,
    output logic [`DATA_WIDTH-1:0]              data_bram_din,
    input  wire [`DATA_WIDTH-1:0]               data_bram_dout
);

    // --- AXI Control Registers ---
    // These will be memory-mapped for the PS to access.
    // Address Map:
    // 0x00 : Control Register (bit 0: start, bit 1: soft_reset)
    // 0x04 : Status Register (bit 0: done)
    // 0x08 : base_instr_addr
    // 0x0C : base_data_addr
    // 0x10 : num_blocks
    // 0x14 : warps_per_block

    logic execution_start_pulse;
    logic soft_reset;
    logic execution_done;

    logic [31:0] base_instr_reg;
    logic [31:0] base_data_reg;
    logic [31:0] num_blocks_reg;
    logic [31:0] warps_per_block_reg;

    // Instantiate the AXI Lite IP generated by Vivado's "Create and Package IP" tool
    // This part is automatically generated by the tool, so we just map the signals.
    // For now, let's create a simple register logic that the real IP will replace.

    wire axi_clk = S_AXI_ACLK;
    wire axi_reset = ~S_AXI_ARESETN;

    // Simple AXI Lite Slave Logic (for simulation, real one generated by Vivado)
    // This logic allows PS to write to our control registers and read status.
    reg_if_axilite #(
        .ADDR_WIDTH(C_S_AXI_ADDR_WIDTH),
        .DATA_WIDTH(C_S_AXI_DATA_WIDTH)
    ) axi_if (
        .clk(axi_clk),
        .reset(axi_reset),
        // AXI signals
        .s_axi_awaddr(S_AXI_AWADDR), .s_axi_awvalid(S_AXI_AWVALID), .s_axi_awready(S_AXI_AWREADY),
        .s_axi_wdata(S_AXI_WDATA), .s_axi_wstrb(S_AXI_WSTRB), .s_axi_wvalid(S_AXI_WVALID), .s_axi_wready(S_AXI_WREADY),
        .s_axi_bresp(S_AXI_BRESP), .s_axi_bvalid(S_AXI_BVALID), .s_axi_bready(S_AXI_BREADY),
        .s_axi_araddr(S_AXI_ARADDR), .s_axi_arvalid(S_AXI_ARVALID), .s_axi_arready(S_AXI_ARREADY),
        .s_axi_rdata(S_AXI_RDATA), .s_axi_rresp(S_AXI_RRESP), .s_axi_rvalid(S_AXI_RVALID), .s_axi_rready(S_AXI_RREADY),
        // Register connections
        .reg0_wdata(S_AXI_WDATA), // Control
        .reg0_rdata({31'b0, execution_done}), // Status
        .reg1_wdata(base_instr_reg),
        .reg1_rdata(base_instr_reg),
        .reg2_wdata(base_data_reg),
        .reg2_rdata(base_data_reg),
        .reg3_wdata(num_blocks_reg),
        .reg3_rdata(num_blocks_reg),
        .reg4_wdata(warps_per_block_reg),
        .reg4_rdata(warps_per_block_reg)
    );
    
    // Create a single-cycle pulse for start
    assign execution_start_pulse = (S_AXI_WVALID && S_AXI_WSTRB[0] && S_AXI_AWADDR == 5'h00 && S_AXI_WDATA[0]);
    assign soft_reset = (S_AXI_WVALID && S_AXI_WSTRB[0] && S_AXI_AWADDR == 5'h00 && S_AXI_WDATA[1]);

    // --- Instantiate GPU and Adapters ---

    // Instruction memory signals
    logic [INSTRUCTION_MEM_NUM_CHANNELS-1:0] imem_valid;
    instruction_memory_address_t imem_addr [INSTRUCTION_MEM_NUM_CHANNELS];
    logic [INSTRUCTION_MEM_NUM_CHANNELS-1:0] imem_ready;
    instruction_t imem_data [INSTRUCTION_MEM_NUM_CHANNELS];

    // Data memory signals
    logic [DATA_MEM_NUM_CHANNELS-1:0] dmem_r_valid;
    data_memory_address_t dmem_r_addr [DATA_MEM_NUM_CHANNELS];
    logic [DATA_MEM_NUM_CHANNELS-1:0] dmem_r_ready;
    data_t dmem_r_data [DATA_MEM_NUM_CHANNELS];
    logic [DATA_MEM_NUM_CHANNELS-1:0] dmem_w_valid;
    data_memory_address_t dmem_w_addr [DATA_MEM_NUM_CHANNELS];
    data_t dmem_w_data [DATA_MEM_NUM_CHANNELS];
    logic [DATA_MEM_NUM_CHANNELS-1:0] dmem_w_ready;


    gpu #(
        .DATA_MEM_NUM_CHANNELS(DATA_MEM_NUM_CHANNELS),
        .INSTRUCTION_MEM_NUM_CHANNELS(INSTRUCTION_MEM_NUM_CHANNELS),
        .NUM_CORES(NUM_CORES),
        .WARPS_PER_CORE(WARPS_PER_CORE),
        .THREADS_PER_WARP(THREADS_PER_WARP)
    ) gpu_inst (
        .clk(axi_clk),
        .reset(axi_reset || soft_reset),
        
        // Kernel Config from AXI regs
        .base_instr(base_instr_reg),
        .base_data(base_data_reg),
        .num_blocks(num_blocks_reg),
        .warps_per_block(warps_per_block_reg),
        
        .execution_start(execution_start_pulse),
        .execution_done(execution_done),

        // Instruction Memory
        .instruction_mem_read_valid(imem_valid),
        .instruction_mem_read_address(imem_addr),
        .instruction_mem_read_ready(imem_ready),
        .instruction_mem_read_data(imem_data),

        // Data Memory
        .data_mem_read_valid(dmem_r_valid),
        .data_mem_read_address(dmem_r_addr),
        .data_mem_read_ready(dmem_r_ready),
        .data_mem_read_data(dmem_r_data),
        .data_mem_write_valid(dmem_w_valid),
        .data_mem_write_address(dmem_w_addr),
        .data_mem_write_data(dmem_w_data),
        .data_mem_write_ready(dmem_w_ready)
    );

    // Adapter for Instruction Memory (Read-Only)
    bram_adapter #(
        .DATA_WIDTH(`INSTRUCTION_WIDTH),
        .ADDR_WIDTH(`INSTRUCTION_MEMORY_ADDRESS_WIDTH),
        .NUM_CHANNELS(INSTRUCTION_MEM_NUM_CHANNELS),
        .WRITE_ENABLE(0)
    ) instr_adapter (
        .clk(axi_clk),
        .reset(axi_reset),
        .gpu_req_valid(imem_valid),
        .gpu_req_ready(imem_ready),
        .gpu_req_addr(imem_addr),
        .gpu_resp_data(imem_data),
        .gpu_w_valid('0), // Not used
        .gpu_w_data('0), // Not used
        .gpu_w_ready(),   // Not used
        .bram_en(instr_bram_en),
        .bram_addr(instr_bram_addr),
        .bram_we(),       // Not used
        .bram_din(),      // Not used
        .bram_dout(instr_bram_dout)
    );

    // Adapter for Data Memory (Read/Write)
    // We combine read and write requests for the arbiter
    logic [DATA_MEM_NUM_CHANNELS-1:0] dmem_any_req_valid;
    data_memory_address_t dmem_any_addr [DATA_MEM_NUM_CHANNELS];
    
    for (genvar i = 0; i < DATA_MEM_NUM_CHANNELS; i++) begin
        assign dmem_any_req_valid[i] = dmem_r_valid[i] || dmem_w_valid[i];
        assign dmem_any_addr[i] = dmem_r_valid[i] ? dmem_r_addr[i] : dmem_w_addr[i];
    end

    bram_adapter #(
        .DATA_WIDTH(`DATA_WIDTH),
        .ADDR_WIDTH(`DATA_MEMORY_ADDRESS_WIDTH),
        .NUM_CHANNELS(DATA_MEM_NUM_CHANNELS),
        .WRITE_ENABLE(1)
    ) data_adapter (
        .clk(axi_clk),
        .reset(axi_reset),
        .gpu_req_valid(dmem_any_req_valid), // Combined read/write valid
        .gpu_req_ready(dmem_r_ready), // Connect ready to both read and write sides
        .gpu_req_addr(dmem_any_addr),
        .gpu_resp_data(dmem_r_data),
        .gpu_w_valid(dmem_w_valid),
        .gpu_w_data(dmem_w_data),
        .gpu_w_ready(dmem_w_ready),
        .bram_en(data_bram_en),
        .bram_addr(data_bram_addr),
        .bram_we(data_bram_we),
        .bram_din(data_bram_din),
        .bram_dout(data_bram_dout)
    );

endmodule

// NOTE: You will need a simple AXI lite slave module like the one that can be generated
// from Vivado's IP templates. For now, this placeholder illustrates the connections.
// To get a real one, use Tools -> Create and Package New IP -> Create AXI4 Peripheral.
`default_nettype wire