module data_mem (
    input  logic                    clk,
    input  logic                    WDME,
    input  logic [31:0]   A,
    input  logic [31:0]   WD,
    output logic [31:0]   RD
);
endmodule